`timescale  1ns/1ns


module  vga_pic
(
    input   wire            vga_clk     ,   //输入工作时钟,频率25MHz
    input   wire            sys_rst_n   ,   //输入复位信号,低电平有效
    input   wire    [9:0]   pix_x       ,   //输入有效显示区域像素点X轴坐标
    input   wire    [9:0]   pix_y       ,   //输入有效显示区域像素点Y轴坐标

    output  reg     [15:0]  pix_data        //输出像素点色彩信息
);


//parameter define
parameter   CHAR_B_H=   10'd192 ,   //字符开始X轴坐标
            CHAR_B_V=   10'd208 ;   //字符开始Y轴坐标

parameter   CHAR_W  =   10'd256 ,   //字符宽度
            CHAR_H  =   10'd64  ;   //字符高度

parameter   BLACK   =   16'h0000,   //黑色
            WHITE   =   16'hFFFF,   //白色
            GOLDEN  =   16'hFEC0;   //金色

//wire  define
wire    [9:0]   char_x  ;   //字符显示X轴坐标
wire    [9:0]   char_y  ;   //字符显示Y轴坐标

//reg   define
reg     [255:0] char    [63:0]  ;   //字符数据



//字符显示坐标
assign  char_x  =   (((pix_x >= CHAR_B_H) && (pix_x < (CHAR_B_H + CHAR_W)))
                    && ((pix_y >= CHAR_B_V) && (pix_y < (CHAR_B_V + CHAR_H))))
                    ? (pix_x - CHAR_B_H) : 10'h3FF;
assign  char_y  =   (((pix_x >= CHAR_B_H) && (pix_x < (CHAR_B_H + CHAR_W)))
                    && ((pix_y >= CHAR_B_V) && (pix_y < (CHAR_B_V + CHAR_H))))
                    ? (pix_y - CHAR_B_V) : 10'h3FF;

//char:字符数据
always@(posedge vga_clk)
    begin
char[0]  <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[1]  <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[2]  <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[3]  <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[4]  <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[5]  <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[6]  <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[7]  <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[8]  <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[9]  <= 256'h00000000000000000000000000000000000003FF000000000000000000000000;
char[10]  <= 256'h7FFC000000FFFE003FFFF80003FFF8000000FFFFFC18000001FFFFFFFFFF8000;
char[11]  <= 256'h03FC000000FFC00001FF0000001F00000007C0007FF8000003FE00FE007F8000;
char[12]  <= 256'h01FE000001FF800000FE0000000E0000001E000007FC000003E000FE000FC000;
char[13]  <= 256'h01FE000001FF800000FE0000000E0000007C000001FC000007C000FE0003C000;
char[14]  <= 256'h01FF000003FF800000FE0000000E000000F8000000FC0000078000FE0001E000;
char[15]  <= 256'h01FF000003BF800000FE0000000E000001F00000007C00000F0000FE0000E000;
char[16]  <= 256'h01BF000003BF800000FE0000000E000003F00000001C00000E0000FE0000E000;
char[17]  <= 256'h019F8000073F800000FE0000000E000003E00000000E00001C0000FE00007000;
char[18]  <= 256'h019F8000073F800000FE0000000E000003E00000000C0000000000FE00000000;
char[19]  <= 256'h018FC0000E3F800000FE0000000E000003F0000000000000000000FE00000000;
char[20]  <= 256'h018FC0000E3F800000FE0000000E000003F0000000000000000000FE00000000;
char[21]  <= 256'h018FE0001C3F800000FE0000000E000003FC000000000000000000FE00000000;
char[22]  <= 256'h0187E0001C3F800000FE0000000E000001FF000000000000000000FE00000000;
char[23]  <= 256'h0187F000383F800000FE0000000E000000FFE00000000000000000FE00000000;
char[24]  <= 256'h0183F000383F800000FE0000000E0000003FFE0000000000000000FE00000000;
char[25]  <= 256'h0183F000703F800000FE0000000E0000000FFFE000000000000000FE00000000;
char[26]  <= 256'h0181F800703F800000FE0000000E00000000FFFE00000000000000FE00000000;
char[27]  <= 256'h0181F800E03F800000FE0000000E000000001FFFF0000000000000FE00000000;
char[28]  <= 256'h0181FC00E03F800000FE0000000E0000000001FFFE000000000000FE00000000;
char[29]  <= 256'h0180FC00E03F800000FE0000000E00000000000FFFC00000000000FE00000000;
char[30]  <= 256'h0180FE01C03F800000FE0000000E000000000000FFF00000000000FE00000000;
char[31]  <= 256'h01807E01C03F800000FE0000000E0000000000001FFC0000000000FE00000000;
char[32]  <= 256'h01807E03803F800000FE0000000E00000000000003FE0000000000FE00000000;
char[33]  <= 256'h01803F03803F800000FE0000000E00000000000000FF0000000000FE00000000;
char[34]  <= 256'h01803F07003F800000FE0000000E000000000000007F8000000000FE00000000;
char[35]  <= 256'h01801F87003F800000FE0000000E000000000000003F8000000000FE00000000;
char[36]  <= 256'h01801F8E003F800000FE0000000E000000000000001F8000000000FE00000000;
char[37]  <= 256'h01801FCE003F800000FE0000000E000007000000001F8000000000FE00000000;
char[38]  <= 256'h01800FDC003F800000FE0000000E000007800000001F8000000000FE00000000;
char[39]  <= 256'h01800FFC003F800000FE0000000E000003C00000001F8000000000FE00000000;
char[40]  <= 256'h018007F8003F800000FE0000000C000003E00000001F8000000000FE00000000;
char[41]  <= 256'h018007F8003F8000007F0000001C000003F00000003F0000000000FE00000000;
char[42]  <= 256'h018003F0003F8000007F00000038000001F80000007E0000000000FE00000000;
char[43]  <= 256'h018003F0003F8000003F800000F0000001FE000000FC0000000000FE00000000;
char[44]  <= 256'h038003E0003F8000000FE00007C0000001FFC00003F00000000000FE00000000;
char[45]  <= 256'h07E001E0007FC0000003FE007F00000000FFFC001FC00000000001FF80000000;
char[46]  <= 256'h7FFC01E00FFFFE0000003FFFF800000000E01FFFFE0000000000FFFFFE000000;
char[47]  <= 256'h00000000000000000000007C000000000000003E000000000000000000000000;
char[48]  <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[49]  <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[50]  <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[51]  <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[52]  <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[53]  <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[54]  <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[55]  <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[56]  <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[57]  <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[58]  <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[59]  <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[60]  <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[61]  <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[62]  <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[63]  <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
end
//pix_data:输出像素点色彩信息,根据当前像素点坐标指定当前像素点颜色数据
always@(posedge vga_clk or negedge sys_rst_n)
    if(sys_rst_n == 1'b0)
        pix_data    <= BLACK;
    else    if((((pix_x >= (CHAR_B_H - 1'b1))
                && (pix_x < (CHAR_B_H + CHAR_W -1'b1)))
                && ((pix_y >= CHAR_B_V) && (pix_y < (CHAR_B_V + CHAR_H))))
                && (char[char_y][10'd255 - char_x] == 1'b1))
        pix_data    <=  GOLDEN;
    else
        pix_data    <=  BLACK;

endmodule
